-- HDMI_QSYS.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HDMI_QSYS is
	port (
		clk_clk                                  : in    std_logic                     := '0'; --                               clk.clk
		hdmi_tx_int_n_external_connection_export : in    std_logic                     := '0'; -- hdmi_tx_int_n_external_connection.export
		i2c_scl_external_connection_export       : out   std_logic;                            --       i2c_scl_external_connection.export
		i2c_sda_external_connection_export       : inout std_logic                     := '0'; --       i2c_sda_external_connection.export
		led_external_connection_export           : out   std_logic_vector(7 downto 0);         --           led_external_connection.export
		position_table_export                    : out   std_logic_vector(31 downto 0);        --                    position_table.export
		refresh_image_export                     : in    std_logic                     := '0'; --                     refresh_image.export
		reset_reset_n                            : in    std_logic                     := '0'  --                             reset.reset_n
	);
end entity HDMI_QSYS;

architecture rtl of HDMI_QSYS is
	component HDMI_QSYS_hdmi_tx_int_n is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component HDMI_QSYS_hdmi_tx_int_n;

	component HDMI_QSYS_i2c_scl is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component HDMI_QSYS_i2c_scl;

	component HDMI_QSYS_i2c_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component HDMI_QSYS_i2c_sda;

	component HDMI_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component HDMI_QSYS_jtag_uart;

	component HDMI_QSYS_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component HDMI_QSYS_led;

	component HDMI_QSYS_nios2_qsys is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(20 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component HDMI_QSYS_nios2_qsys;

	component HDMI_QSYS_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component HDMI_QSYS_onchip_memory2;

	component HDMI_QSYS_pll_sys is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component HDMI_QSYS_pll_sys;

	component HDMI_QSYS_position is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component HDMI_QSYS_position;

	component HDMI_QSYS_refresh is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component HDMI_QSYS_refresh;

	component HDMI_QSYS_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component HDMI_QSYS_sysid_qsys;

	component HDMI_QSYS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component HDMI_QSYS_timer;

	component HDMI_QSYS_mm_interconnect_0 is
		port (
			clk_50_clk_clk                               : in  std_logic                     := 'X';             -- clk
			pll_sys_outclk0_clk                          : in  std_logic                     := 'X';             -- clk
			nios2_qsys_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			position_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			nios2_qsys_data_master_address               : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_qsys_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_qsys_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_qsys_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_qsys_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_qsys_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_instruction_master_address        : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_qsys_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_qsys_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_qsys_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			hdmi_tx_int_n_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			hdmi_tx_int_n_s1_write                       : out std_logic;                                        -- write
			hdmi_tx_int_n_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hdmi_tx_int_n_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			hdmi_tx_int_n_s1_chipselect                  : out std_logic;                                        -- chipselect
			i2c_scl_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			i2c_scl_s1_write                             : out std_logic;                                        -- write
			i2c_scl_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_scl_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_scl_s1_chipselect                        : out std_logic;                                        -- chipselect
			i2c_sda_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			i2c_sda_s1_write                             : out std_logic;                                        -- write
			i2c_sda_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_sda_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_sda_s1_chipselect                        : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			led_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                 : out std_logic;                                        -- write
			led_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                            : out std_logic;                                        -- chipselect
			nios2_qsys_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_qsys_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_qsys_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_s1_address                    : out std_logic_vector(16 downto 0);                    -- address
			onchip_memory2_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                      : out std_logic;                                        -- clken
			position_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			position_s1_write                            : out std_logic;                                        -- write
			position_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			position_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			position_s1_chipselect                       : out std_logic;                                        -- chipselect
			refresh_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			refresh_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                             : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                               : out std_logic;                                        -- write
			timer_s1_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                          : out std_logic                                         -- chipselect
		);
	end component HDMI_QSYS_mm_interconnect_0;

	component HDMI_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component HDMI_QSYS_irq_mapper;

	component hdmi_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component hdmi_qsys_rst_controller;

	component hdmi_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component hdmi_qsys_rst_controller_001;

	signal pll_sys_outclk0_clk                                           : std_logic;                     -- pll_sys:outclk_0 -> [hdmi_tx_int_n:clk, i2c_scl:clk, i2c_sda:clk, irq_mapper:clk, jtag_uart:clk, led:clk, mm_interconnect_0:pll_sys_outclk0_clk, nios2_qsys:clk, onchip_memory2:clk, rst_controller:clk, sysid_qsys:clock, timer:clk]
	signal nios2_qsys_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_debugaccess                            : std_logic;                     -- nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	signal nios2_qsys_data_master_address                                : std_logic_vector(20 downto 0); -- nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	signal nios2_qsys_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	signal nios2_qsys_data_master_read                                   : std_logic;                     -- nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	signal nios2_qsys_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	signal nios2_qsys_data_master_write                                  : std_logic;                     -- nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	signal nios2_qsys_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	signal nios2_qsys_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                         : std_logic_vector(20 downto 0); -- nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	signal nios2_qsys_instruction_master_read                            : std_logic;                     -- nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	signal nios2_qsys_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                   : std_logic_vector(16 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_i2c_sda_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	signal mm_interconnect_0_i2c_sda_s1_readdata                         : std_logic_vector(31 downto 0); -- i2c_sda:readdata -> mm_interconnect_0:i2c_sda_s1_readdata
	signal mm_interconnect_0_i2c_sda_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:i2c_sda_s1_address -> i2c_sda:address
	signal mm_interconnect_0_i2c_sda_s1_write                            : std_logic;                     -- mm_interconnect_0:i2c_sda_s1_write -> mm_interconnect_0_i2c_sda_s1_write:in
	signal mm_interconnect_0_i2c_sda_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:i2c_sda_s1_writedata -> i2c_sda:writedata
	signal mm_interconnect_0_i2c_scl_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	signal mm_interconnect_0_i2c_scl_s1_readdata                         : std_logic_vector(31 downto 0); -- i2c_scl:readdata -> mm_interconnect_0:i2c_scl_s1_readdata
	signal mm_interconnect_0_i2c_scl_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:i2c_scl_s1_address -> i2c_scl:address
	signal mm_interconnect_0_i2c_scl_s1_write                            : std_logic;                     -- mm_interconnect_0:i2c_scl_s1_write -> mm_interconnect_0_i2c_scl_s1_write:in
	signal mm_interconnect_0_i2c_scl_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:i2c_scl_s1_writedata -> i2c_scl:writedata
	signal mm_interconnect_0_led_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                             : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_hdmi_tx_int_n_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:hdmi_tx_int_n_s1_chipselect -> hdmi_tx_int_n:chipselect
	signal mm_interconnect_0_hdmi_tx_int_n_s1_readdata                   : std_logic_vector(31 downto 0); -- hdmi_tx_int_n:readdata -> mm_interconnect_0:hdmi_tx_int_n_s1_readdata
	signal mm_interconnect_0_hdmi_tx_int_n_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hdmi_tx_int_n_s1_address -> hdmi_tx_int_n:address
	signal mm_interconnect_0_hdmi_tx_int_n_s1_write                      : std_logic;                     -- mm_interconnect_0:hdmi_tx_int_n_s1_write -> mm_interconnect_0_hdmi_tx_int_n_s1_write:in
	signal mm_interconnect_0_hdmi_tx_int_n_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hdmi_tx_int_n_s1_writedata -> hdmi_tx_int_n:writedata
	signal mm_interconnect_0_position_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:position_s1_chipselect -> position:chipselect
	signal mm_interconnect_0_position_s1_readdata                        : std_logic_vector(31 downto 0); -- position:readdata -> mm_interconnect_0:position_s1_readdata
	signal mm_interconnect_0_position_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:position_s1_address -> position:address
	signal mm_interconnect_0_position_s1_write                           : std_logic;                     -- mm_interconnect_0:position_s1_write -> mm_interconnect_0_position_s1_write:in
	signal mm_interconnect_0_position_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:position_s1_writedata -> position:writedata
	signal mm_interconnect_0_refresh_s1_readdata                         : std_logic_vector(31 downto 0); -- refresh:readdata -> mm_interconnect_0:refresh_s1_readdata
	signal mm_interconnect_0_refresh_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:refresh_s1_address -> refresh:address
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- timer:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- hdmi_tx_int_n:irq -> irq_mapper:receiver2_irq
	signal nios2_qsys_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [nios2_qsys:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:position_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [pll_sys:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_0_i2c_sda_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_i2c_sda_s1_write:inv -> i2c_sda:write_n
	signal mm_interconnect_0_i2c_scl_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_i2c_scl_s1_write:inv -> i2c_scl:write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_hdmi_tx_int_n_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_hdmi_tx_int_n_s1_write:inv -> hdmi_tx_int_n:write_n
	signal mm_interconnect_0_position_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_position_s1_write:inv -> position:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [hdmi_tx_int_n:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, jtag_uart:rst_n, led:reset_n, nios2_qsys:reset_n, sysid_qsys:reset_n, timer:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [position:reset_n, refresh:reset_n]

begin

	hdmi_tx_int_n : component HDMI_QSYS_hdmi_tx_int_n
		port map (
			clk        => pll_sys_outclk0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_hdmi_tx_int_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hdmi_tx_int_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hdmi_tx_int_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hdmi_tx_int_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hdmi_tx_int_n_s1_readdata,        --                    .readdata
			in_port    => hdmi_tx_int_n_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                            --                 irq.irq
		);

	i2c_scl : component HDMI_QSYS_i2c_scl
		port map (
			clk        => pll_sys_outclk0_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => i2c_scl_external_connection_export            -- external_connection.export
		);

	i2c_sda : component HDMI_QSYS_i2c_sda
		port map (
			clk        => pll_sys_outclk0_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => i2c_sda_external_connection_export            -- external_connection.export
		);

	jtag_uart : component HDMI_QSYS_jtag_uart
		port map (
			clk            => pll_sys_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	led : component HDMI_QSYS_led
		port map (
			clk        => pll_sys_outclk0_clk,                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	nios2_qsys : component HDMI_QSYS_nios2_qsys
		port map (
			clk                                 => pll_sys_outclk0_clk,                                      --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
			d_address                           => nios2_qsys_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_qsys_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_qsys_data_master_read,                              --                          .read
			d_readdata                          => nios2_qsys_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_qsys_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_qsys_data_master_write,                             --                          .write
			d_writedata                         => nios2_qsys_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_qsys_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_qsys_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_qsys_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_qsys_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_qsys_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_qsys_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_qsys_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_qsys_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_qsys_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_qsys_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	onchip_memory2 : component HDMI_QSYS_onchip_memory2
		port map (
			clk        => pll_sys_outclk0_clk,                            --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	pll_sys : component HDMI_QSYS_pll_sys
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_sys_outclk0_clk,     -- outclk0.clk
			locked   => open                     --  locked.export
		);

	position : component HDMI_QSYS_position
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_position_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_position_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_position_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_position_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_position_s1_readdata,        --                    .readdata
			out_port   => position_table_export                          -- external_connection.export
		);

	refresh : component HDMI_QSYS_refresh
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_refresh_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_refresh_s1_readdata,        --                    .readdata
			in_port  => refresh_image_export                          -- external_connection.export
		);

	sysid_qsys : component HDMI_QSYS_sysid_qsys
		port map (
			clock    => pll_sys_outclk0_clk,                                   --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer : component HDMI_QSYS_timer
		port map (
			clk        => pll_sys_outclk0_clk,                        --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                    --   irq.irq
		);

	mm_interconnect_0 : component HDMI_QSYS_mm_interconnect_0
		port map (
			clk_50_clk_clk                               => clk_clk,                                                   --                             clk_50_clk.clk
			pll_sys_outclk0_clk                          => pll_sys_outclk0_clk,                                       --                        pll_sys_outclk0.clk
			nios2_qsys_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- nios2_qsys_reset_reset_bridge_in_reset.reset
			position_reset_reset_bridge_in_reset_reset   => rst_controller_001_reset_out_reset,                        --   position_reset_reset_bridge_in_reset.reset
			nios2_qsys_data_master_address               => nios2_qsys_data_master_address,                            --                 nios2_qsys_data_master.address
			nios2_qsys_data_master_waitrequest           => nios2_qsys_data_master_waitrequest,                        --                                       .waitrequest
			nios2_qsys_data_master_byteenable            => nios2_qsys_data_master_byteenable,                         --                                       .byteenable
			nios2_qsys_data_master_read                  => nios2_qsys_data_master_read,                               --                                       .read
			nios2_qsys_data_master_readdata              => nios2_qsys_data_master_readdata,                           --                                       .readdata
			nios2_qsys_data_master_readdatavalid         => nios2_qsys_data_master_readdatavalid,                      --                                       .readdatavalid
			nios2_qsys_data_master_write                 => nios2_qsys_data_master_write,                              --                                       .write
			nios2_qsys_data_master_writedata             => nios2_qsys_data_master_writedata,                          --                                       .writedata
			nios2_qsys_data_master_debugaccess           => nios2_qsys_data_master_debugaccess,                        --                                       .debugaccess
			nios2_qsys_instruction_master_address        => nios2_qsys_instruction_master_address,                     --          nios2_qsys_instruction_master.address
			nios2_qsys_instruction_master_waitrequest    => nios2_qsys_instruction_master_waitrequest,                 --                                       .waitrequest
			nios2_qsys_instruction_master_read           => nios2_qsys_instruction_master_read,                        --                                       .read
			nios2_qsys_instruction_master_readdata       => nios2_qsys_instruction_master_readdata,                    --                                       .readdata
			nios2_qsys_instruction_master_readdatavalid  => nios2_qsys_instruction_master_readdatavalid,               --                                       .readdatavalid
			hdmi_tx_int_n_s1_address                     => mm_interconnect_0_hdmi_tx_int_n_s1_address,                --                       hdmi_tx_int_n_s1.address
			hdmi_tx_int_n_s1_write                       => mm_interconnect_0_hdmi_tx_int_n_s1_write,                  --                                       .write
			hdmi_tx_int_n_s1_readdata                    => mm_interconnect_0_hdmi_tx_int_n_s1_readdata,               --                                       .readdata
			hdmi_tx_int_n_s1_writedata                   => mm_interconnect_0_hdmi_tx_int_n_s1_writedata,              --                                       .writedata
			hdmi_tx_int_n_s1_chipselect                  => mm_interconnect_0_hdmi_tx_int_n_s1_chipselect,             --                                       .chipselect
			i2c_scl_s1_address                           => mm_interconnect_0_i2c_scl_s1_address,                      --                             i2c_scl_s1.address
			i2c_scl_s1_write                             => mm_interconnect_0_i2c_scl_s1_write,                        --                                       .write
			i2c_scl_s1_readdata                          => mm_interconnect_0_i2c_scl_s1_readdata,                     --                                       .readdata
			i2c_scl_s1_writedata                         => mm_interconnect_0_i2c_scl_s1_writedata,                    --                                       .writedata
			i2c_scl_s1_chipselect                        => mm_interconnect_0_i2c_scl_s1_chipselect,                   --                                       .chipselect
			i2c_sda_s1_address                           => mm_interconnect_0_i2c_sda_s1_address,                      --                             i2c_sda_s1.address
			i2c_sda_s1_write                             => mm_interconnect_0_i2c_sda_s1_write,                        --                                       .write
			i2c_sda_s1_readdata                          => mm_interconnect_0_i2c_sda_s1_readdata,                     --                                       .readdata
			i2c_sda_s1_writedata                         => mm_interconnect_0_i2c_sda_s1_writedata,                    --                                       .writedata
			i2c_sda_s1_chipselect                        => mm_interconnect_0_i2c_sda_s1_chipselect,                   --                                       .chipselect
			jtag_uart_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --            jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                       .write
			jtag_uart_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                       .read
			jtag_uart_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                       .readdata
			jtag_uart_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                       .writedata
			jtag_uart_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                       .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                       .chipselect
			led_s1_address                               => mm_interconnect_0_led_s1_address,                          --                                 led_s1.address
			led_s1_write                                 => mm_interconnect_0_led_s1_write,                            --                                       .write
			led_s1_readdata                              => mm_interconnect_0_led_s1_readdata,                         --                                       .readdata
			led_s1_writedata                             => mm_interconnect_0_led_s1_writedata,                        --                                       .writedata
			led_s1_chipselect                            => mm_interconnect_0_led_s1_chipselect,                       --                                       .chipselect
			nios2_qsys_debug_mem_slave_address           => mm_interconnect_0_nios2_qsys_debug_mem_slave_address,      --             nios2_qsys_debug_mem_slave.address
			nios2_qsys_debug_mem_slave_write             => mm_interconnect_0_nios2_qsys_debug_mem_slave_write,        --                                       .write
			nios2_qsys_debug_mem_slave_read              => mm_interconnect_0_nios2_qsys_debug_mem_slave_read,         --                                       .read
			nios2_qsys_debug_mem_slave_readdata          => mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata,     --                                       .readdata
			nios2_qsys_debug_mem_slave_writedata         => mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata,    --                                       .writedata
			nios2_qsys_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable,   --                                       .byteenable
			nios2_qsys_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest,  --                                       .waitrequest
			nios2_qsys_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess,  --                                       .debugaccess
			onchip_memory2_s1_address                    => mm_interconnect_0_onchip_memory2_s1_address,               --                      onchip_memory2_s1.address
			onchip_memory2_s1_write                      => mm_interconnect_0_onchip_memory2_s1_write,                 --                                       .write
			onchip_memory2_s1_readdata                   => mm_interconnect_0_onchip_memory2_s1_readdata,              --                                       .readdata
			onchip_memory2_s1_writedata                  => mm_interconnect_0_onchip_memory2_s1_writedata,             --                                       .writedata
			onchip_memory2_s1_byteenable                 => mm_interconnect_0_onchip_memory2_s1_byteenable,            --                                       .byteenable
			onchip_memory2_s1_chipselect                 => mm_interconnect_0_onchip_memory2_s1_chipselect,            --                                       .chipselect
			onchip_memory2_s1_clken                      => mm_interconnect_0_onchip_memory2_s1_clken,                 --                                       .clken
			position_s1_address                          => mm_interconnect_0_position_s1_address,                     --                            position_s1.address
			position_s1_write                            => mm_interconnect_0_position_s1_write,                       --                                       .write
			position_s1_readdata                         => mm_interconnect_0_position_s1_readdata,                    --                                       .readdata
			position_s1_writedata                        => mm_interconnect_0_position_s1_writedata,                   --                                       .writedata
			position_s1_chipselect                       => mm_interconnect_0_position_s1_chipselect,                  --                                       .chipselect
			refresh_s1_address                           => mm_interconnect_0_refresh_s1_address,                      --                             refresh_s1.address
			refresh_s1_readdata                          => mm_interconnect_0_refresh_s1_readdata,                     --                                       .readdata
			sysid_qsys_control_slave_address             => mm_interconnect_0_sysid_qsys_control_slave_address,        --               sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata            => mm_interconnect_0_sysid_qsys_control_slave_readdata,       --                                       .readdata
			timer_s1_address                             => mm_interconnect_0_timer_s1_address,                        --                               timer_s1.address
			timer_s1_write                               => mm_interconnect_0_timer_s1_write,                          --                                       .write
			timer_s1_readdata                            => mm_interconnect_0_timer_s1_readdata,                       --                                       .readdata
			timer_s1_writedata                           => mm_interconnect_0_timer_s1_writedata,                      --                                       .writedata
			timer_s1_chipselect                          => mm_interconnect_0_timer_s1_chipselect                      --                                       .chipselect
		);

	irq_mapper : component HDMI_QSYS_irq_mapper
		port map (
			clk           => pll_sys_outclk0_clk,            --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_qsys_irq_irq              --    sender.irq
		);

	rst_controller : component hdmi_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_sys_outclk0_clk,                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component hdmi_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_i2c_sda_s1_write_ports_inv <= not mm_interconnect_0_i2c_sda_s1_write;

	mm_interconnect_0_i2c_scl_s1_write_ports_inv <= not mm_interconnect_0_i2c_scl_s1_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_hdmi_tx_int_n_s1_write_ports_inv <= not mm_interconnect_0_hdmi_tx_int_n_s1_write;

	mm_interconnect_0_position_s1_write_ports_inv <= not mm_interconnect_0_position_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of HDMI_QSYS
