-- nios_arch.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_arch is
	port (
		nios2_qsys_0_custom_instruction_master_readra : out   std_logic;                                        -- nios2_qsys_0_custom_instruction_master.readra
		nios2_qsys_0_d_irq_irq                        : in    std_logic_vector(31 downto 0) := (others => '0'); --                     nios2_qsys_0_d_irq.irq
		terasic_sram_0_conduit_end_DQ                 : inout std_logic_vector(15 downto 0) := (others => '0'); --             terasic_sram_0_conduit_end.DQ
		terasic_sram_0_conduit_end_ADDR               : out   std_logic_vector(19 downto 0);                    --                                       .ADDR
		terasic_sram_0_conduit_end_UB_n               : out   std_logic;                                        --                                       .UB_n
		terasic_sram_0_conduit_end_LB_n               : out   std_logic;                                        --                                       .LB_n
		terasic_sram_0_conduit_end_WE_n               : out   std_logic;                                        --                                       .WE_n
		terasic_sram_0_conduit_end_CE_n               : out   std_logic;                                        --                                       .CE_n
		terasic_sram_0_conduit_end_OE_n               : out   std_logic                                         --                                       .OE_n
	);
end entity nios_arch;

architecture rtl of nios_arch is
	component TERASIC_SRAM is
		generic (
			DATA_BITS : integer := 16;
			ADDR_BITS : integer := 20
		);
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			s_chipselect_n : in    std_logic                     := 'X';             -- chipselect_n
			s_write_n      : in    std_logic                     := 'X';             -- write_n
			s_address      : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			s_read_n       : in    std_logic                     := 'X';             -- read_n
			s_writedata    : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			s_readdata     : out   std_logic_vector(15 downto 0);                    -- readdata
			s_byteenable_n : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			SRAM_DQ        : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR      : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_UB_n      : out   std_logic;                                        -- export
			SRAM_LB_n      : out   std_logic;                                        -- export
			SRAM_WE_n      : out   std_logic;                                        -- export
			SRAM_CE_n      : out   std_logic;                                        -- export
			SRAM_OE_n      : out   std_logic                                         -- export
		);
	end component TERASIC_SRAM;

	component nios_arch_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(21 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(21 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_arch_nios2_qsys_0;

	component nios_arch_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_arch_onchip_memory2_0;

	component nios_arch_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_data_master_address                 : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address          : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                      : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                        : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                        : out std_logic;                                        -- clken
			TERASIC_SRAM_0_avalon_slave_address              : out std_logic_vector(19 downto 0);                    -- address
			TERASIC_SRAM_0_avalon_slave_write                : out std_logic;                                        -- write
			TERASIC_SRAM_0_avalon_slave_read                 : out std_logic;                                        -- read
			TERASIC_SRAM_0_avalon_slave_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TERASIC_SRAM_0_avalon_slave_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			TERASIC_SRAM_0_avalon_slave_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			TERASIC_SRAM_0_avalon_slave_chipselect           : out std_logic                                         -- chipselect
		);
	end component nios_arch_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal terasic_sram_0_clock_reset_clk                                     : std_logic;                     -- [] -> [TERASIC_SRAM_0:clk, mm_interconnect_0:clk_0_clk_clk, nios2_qsys_0:clk, onchip_memory2_0:clk, rst_controller:clk]
	signal nios2_qsys_0_jtag_debug_module_reset_reset                         : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal nios2_qsys_0_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_debugaccess                               : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_address                                   : std_logic_vector(21 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_data_master_read                                      : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_write                                     : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_writedata                                 : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                            : std_logic_vector(21 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                               : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect           : std_logic;                     -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_chipselect -> mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect:in
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_readdata             : std_logic_vector(15 downto 0); -- TERASIC_SRAM_0:s_readdata -> mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_readdata
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_address              : std_logic_vector(19 downto 0); -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_address -> TERASIC_SRAM_0:s_address
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_read                 : std_logic;                     -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_read -> mm_interconnect_0_terasic_sram_0_avalon_slave_read:in
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_byteenable -> mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable:in
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_write                : std_logic;                     -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_write -> mm_interconnect_0_terasic_sram_0_avalon_slave_write:in
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:TERASIC_SRAM_0_avalon_slave_writedata -> TERASIC_SRAM_0:s_writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata          : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest       : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess       : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read              : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write             : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                     : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                      : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in]
	signal rst_controller_reset_out_reset_req                                 : std_logic;                     -- rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect:inv -> TERASIC_SRAM_0:s_chipselect_n
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_terasic_sram_0_avalon_slave_read:inv -> TERASIC_SRAM_0:s_read_n
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable_ports_inv : std_logic_vector(1 downto 0);  -- mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable:inv -> TERASIC_SRAM_0:s_byteenable_n
	signal mm_interconnect_0_terasic_sram_0_avalon_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_terasic_sram_0_avalon_slave_write:inv -> TERASIC_SRAM_0:s_write_n
	signal rst_controller_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [TERASIC_SRAM_0:reset_n, nios2_qsys_0:reset_n]

begin

	terasic_sram_0 : component TERASIC_SRAM
		generic map (
			DATA_BITS => 16,
			ADDR_BITS => 20
		)
		port map (
			clk            => terasic_sram_0_clock_reset_clk,                                     --       clock_reset.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                           -- clock_reset_reset.reset_n
			s_chipselect_n => mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect_ports_inv, --      avalon_slave.chipselect_n
			s_write_n      => mm_interconnect_0_terasic_sram_0_avalon_slave_write_ports_inv,      --                  .write_n
			s_address      => mm_interconnect_0_terasic_sram_0_avalon_slave_address,              --                  .address
			s_read_n       => mm_interconnect_0_terasic_sram_0_avalon_slave_read_ports_inv,       --                  .read_n
			s_writedata    => mm_interconnect_0_terasic_sram_0_avalon_slave_writedata,            --                  .writedata
			s_readdata     => mm_interconnect_0_terasic_sram_0_avalon_slave_readdata,             --                  .readdata
			s_byteenable_n => mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable_ports_inv, --                  .byteenable_n
			SRAM_DQ        => terasic_sram_0_conduit_end_DQ,                                      --       conduit_end.export
			SRAM_ADDR      => terasic_sram_0_conduit_end_ADDR,                                    --                  .export
			SRAM_UB_n      => terasic_sram_0_conduit_end_UB_n,                                    --                  .export
			SRAM_LB_n      => terasic_sram_0_conduit_end_LB_n,                                    --                  .export
			SRAM_WE_n      => terasic_sram_0_conduit_end_WE_n,                                    --                  .export
			SRAM_CE_n      => terasic_sram_0_conduit_end_CE_n,                                    --                  .export
			SRAM_OE_n      => terasic_sram_0_conduit_end_OE_n                                     --                  .export
		);

	nios2_qsys_0 : component nios_arch_nios2_qsys_0
		port map (
			clk                                   => terasic_sram_0_clock_reset_clk,                               --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                     --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                           --                          .reset_req
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => nios2_qsys_0_custom_instruction_master_readra                 -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component nios_arch_onchip_memory2_0
		port map (
			clk        => terasic_sram_0_clock_reset_clk,                   --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	mm_interconnect_0 : component nios_arch_mm_interconnect_0
		port map (
			clk_0_clk_clk                                    => terasic_sram_0_clock_reset_clk,                               --                                  clk_0_clk.clk
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                               -- nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_0_data_master_address                 => nios2_qsys_0_data_master_address,                             --                   nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest             => nios2_qsys_0_data_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_0_data_master_byteenable              => nios2_qsys_0_data_master_byteenable,                          --                                           .byteenable
			nios2_qsys_0_data_master_read                    => nios2_qsys_0_data_master_read,                                --                                           .read
			nios2_qsys_0_data_master_readdata                => nios2_qsys_0_data_master_readdata,                            --                                           .readdata
			nios2_qsys_0_data_master_write                   => nios2_qsys_0_data_master_write,                               --                                           .write
			nios2_qsys_0_data_master_writedata               => nios2_qsys_0_data_master_writedata,                           --                                           .writedata
			nios2_qsys_0_data_master_debugaccess             => nios2_qsys_0_data_master_debugaccess,                         --                                           .debugaccess
			nios2_qsys_0_instruction_master_address          => nios2_qsys_0_instruction_master_address,                      --            nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest      => nios2_qsys_0_instruction_master_waitrequest,                  --                                           .waitrequest
			nios2_qsys_0_instruction_master_read             => nios2_qsys_0_instruction_master_read,                         --                                           .read
			nios2_qsys_0_instruction_master_readdata         => nios2_qsys_0_instruction_master_readdata,                     --                                           .readdata
			nios2_qsys_0_jtag_debug_module_address           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --             nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                                           .write
			nios2_qsys_0_jtag_debug_module_read              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                                           .read
			nios2_qsys_0_jtag_debug_module_readdata          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                                           .readdata
			nios2_qsys_0_jtag_debug_module_writedata         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                                           .writedata
			nios2_qsys_0_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                                           .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                                           .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                                           .debugaccess
			onchip_memory2_0_s1_address                      => mm_interconnect_0_onchip_memory2_0_s1_address,                --                        onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                        => mm_interconnect_0_onchip_memory2_0_s1_write,                  --                                           .write
			onchip_memory2_0_s1_readdata                     => mm_interconnect_0_onchip_memory2_0_s1_readdata,               --                                           .readdata
			onchip_memory2_0_s1_writedata                    => mm_interconnect_0_onchip_memory2_0_s1_writedata,              --                                           .writedata
			onchip_memory2_0_s1_byteenable                   => mm_interconnect_0_onchip_memory2_0_s1_byteenable,             --                                           .byteenable
			onchip_memory2_0_s1_chipselect                   => mm_interconnect_0_onchip_memory2_0_s1_chipselect,             --                                           .chipselect
			onchip_memory2_0_s1_clken                        => mm_interconnect_0_onchip_memory2_0_s1_clken,                  --                                           .clken
			TERASIC_SRAM_0_avalon_slave_address              => mm_interconnect_0_terasic_sram_0_avalon_slave_address,        --                TERASIC_SRAM_0_avalon_slave.address
			TERASIC_SRAM_0_avalon_slave_write                => mm_interconnect_0_terasic_sram_0_avalon_slave_write,          --                                           .write
			TERASIC_SRAM_0_avalon_slave_read                 => mm_interconnect_0_terasic_sram_0_avalon_slave_read,           --                                           .read
			TERASIC_SRAM_0_avalon_slave_readdata             => mm_interconnect_0_terasic_sram_0_avalon_slave_readdata,       --                                           .readdata
			TERASIC_SRAM_0_avalon_slave_writedata            => mm_interconnect_0_terasic_sram_0_avalon_slave_writedata,      --                                           .writedata
			TERASIC_SRAM_0_avalon_slave_byteenable           => mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable,     --                                           .byteenable
			TERASIC_SRAM_0_avalon_slave_chipselect           => mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect      --                                           .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => terasic_sram_0_clock_reset_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,         --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect_ports_inv <= not mm_interconnect_0_terasic_sram_0_avalon_slave_chipselect;

	mm_interconnect_0_terasic_sram_0_avalon_slave_read_ports_inv <= not mm_interconnect_0_terasic_sram_0_avalon_slave_read;

	mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable_ports_inv <= not mm_interconnect_0_terasic_sram_0_avalon_slave_byteenable;

	mm_interconnect_0_terasic_sram_0_avalon_slave_write_ports_inv <= not mm_interconnect_0_terasic_sram_0_avalon_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_arch
